package count_pkg;  

import uvm_pkg::*;
`include "uvm_macros.svh"
   //`include the files 
`include "count_trans.sv"
`include "count_config.sv"
 `include "count_driver.sv"
 `include "count_monitor.sv"
`include "count_sequencer.sv"
`include "count_agent.sv" 
 `include "count_sb.sv"
 `include "counter_env.sv"
`include "count_seq.sv"
 `include "test.sv" 
endpackage
